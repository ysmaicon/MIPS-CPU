module Register(
	input clock,
	input [31:0] entrada,
	output reg [31:0] saida
	);

	always @(posedge clock)begin
		saida <= entrada;
	end
	
endmodule
